--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   13:41:45 06/16/2020
-- Design Name:   
-- Module Name:   C:/LUCIANO/TESIS/ADS8694_Handler/ADS8694_Handler/ADS8694_Handler/test/fixed_test.vhd
-- Project Name:  ADS8694_Handler
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: SOS
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
library std;
use std.textio.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE ieee.numeric_std.ALL;
 
ENTITY fixed_test IS
END fixed_test;
 
ARCHITECTURE behavior OF fixed_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT SOS
	 	 generic(
		b0	:	signed(31 downto 0) := "00100000000000000000000000000000";
		b1	:	signed(31 downto 0) := "01000000000000000000000000000000";
		b2	:	signed(31 downto 0) := "00100000000000000000000000000000";
		a1	:	signed(31 downto 0) := "11000000001000101011101011011111";
		a2	:	signed(31 downto 0) := "00011111110111100011000001001001";
		g	:	signed(31 downto 0) := "00000000000000000011101011001010"
	 );
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         data_i : IN  std_logic_vector(17 downto 0);
         data_o : OUT  std_logic_vector(18 downto 0);
         data_o_en : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal data_i_1 : std_logic_vector(17 downto 0) := (others => '0');
   signal data_i_2 : std_logic_vector(17 downto 0) := (others => '0');
   signal data_i_3 : std_logic_vector(17 downto 0) := (others => '0');
   signal data_i_4 : std_logic_vector(17 downto 0) := (others => '0');

 	--Outputs
   signal data_o_1 : std_logic_vector(18 downto 0);
   signal data_o_en_1 : std_logic;
   signal data_o_2 : std_logic_vector(18 downto 0);
   signal data_o_en_2 : std_logic;
   signal data_o_3 : std_logic_vector(18 downto 0);
   signal data_o_en_3 : std_logic;
   signal data_o_4 : std_logic_vector(18 downto 0);
   signal data_o_en_4 : std_logic;
		
   -- Clock period definitions
   constant clk_period : time := 50 us;
 
   file f : text;
 
BEGIN
--SOS Matrix:                                                                                                                                                                                               
--00100000000000000000000000000000  01000000000000000000000000000000  00100000000000000000000000000000  00100000000000000000000000000000  11000000001000101011101011011111  00011111110111100011000001001001
--00100000000000000000000000000000  01000000000000000000000000000000  00100000000000000000000000000000  00100000000000000000000000000000  11000000011000001101011000000100  00011111101000000001010000111111
--00100000000000000000000000000000  01000000000000000000000000000000  00100000000000000000000000000000  00100000000000000000000000000000  11000000100100000000110101010100  00011111011100001101110001000001
--00100000000000000000000000000000  01000000000000000000000000000000  00100000000000000000000000000000  00100000000000000000000000000000  11000000101010010111110111000001  00011111010101110110101101110110
--                                                                                                                                                                                                          
--Scale Values:                                                                                                                                                                                             
--00000000000000000011101011001010                                                                                                                                                                          
--00000000000000000011101010010001                                                                                                                                                                          
--00000000000000000011101001100101                                                                                                                                                                          
--00000000000000000011101001001110 
 
	-- Instantiate the Unit Under Test (UUT)
   SOS1: SOS 
	GENERIC MAP(
		b0	=> "00100000000000000000000000000000",
		b1	=> "01000000000000000000000000000000",
		b2	=> "00100000000000000000000000000000",
		a1	=> "11000000001000101011101011011111",
		a2	=> "00011111110111100011000001001001",
		g	=> "00000000000000000011101011001010"
	)
	PORT MAP (
          clk => clk,
          reset => reset,
          data_i => data_i_1,
          data_o => data_o_1,
          data_o_en => data_o_en_1
        );
		  
	SOS2: SOS 
	GENERIC MAP(
		b0	=> "00100000000000000000000000000000",
		b1	=> "01000000000000000000000000000000",
		b2	=> "00100000000000000000000000000000",
		a1	=> "11000000011000001101011000000100",
		a2	=> "00011111101000000001010000111111",
		g	=> "00000000000000000011101010010001"
	)
	PORT MAP (
          clk => clk,
          reset => reset,
          data_i => data_i_2,
          data_o => data_o_2,
          data_o_en => data_o_en_2
        );
		  
		  
	SOS3: SOS 
	GENERIC MAP(
		b0	=> "00100000000000000000000000000000",
		b1	=> "01000000000000000000000000000000",
		b2	=> "00100000000000000000000000000000",
		a1	=> "11000000100100000000110101010100",
		a2	=> "00011111011100001101110001000001",
		g	=> "00000000000000000011101001100101"
	)
	PORT MAP (
          clk => clk,
          reset => reset,
          data_i => data_i_3,
          data_o => data_o_3,
          data_o_en => data_o_en_3
        );
		  
		  
		  
	SOS4: SOS 
	GENERIC MAP(
		b0	=> "00100000000000000000000000000000",
		b1	=> "01000000000000000000000000000000",
		b2	=> "00100000000000000000000000000000",
		a1	=> "11000000101010010111110111000001",
		a2	=> "00011111010101110110101101110110",
		g	=> "00000000000000000011101001001110"
	)
	PORT MAP (
          clk => clk,
          reset => reset,
          data_i => data_i_4,
          data_o => data_o_4,
          data_o_en => data_o_en_4
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

	data_i_2 <= data_o_1(17 downto 0); 
	data_i_3 <= data_o_2(17 downto 0);
	data_i_4 <= data_o_3(17 downto 0);

   -- Stimulus process
   stim_proc: process
		variable l      : line;
      variable status : file_open_status;
	begin
		file_open(status,f,"resul_iir.m",write_mode);
		assert status=open_ok
		report "No se pudo crear resul_iir.m"
		severity failure;
      -- hold reset state for 100 ns.
		reset <= '1';
      wait for clk_period;
		reset <= '0';
		wait until rising_edge(clk);
		wait for clk_period/2;
		wait for clk_period/2;


		
		data_i_1 <= std_logic_vector(to_unsigned(131072,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(133130,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(135189,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(137246,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(139302,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(141355,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(143406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(145455,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(147499,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(149540,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(151576,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(153607,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(155632,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(157651,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(159664,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(161670,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(163668,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(165658,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(167639,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(169612,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(171575,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(173528,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(175470,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(177402,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(179322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(181230,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(183126,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(185009,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(186879,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(188735,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(190577,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(192404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(194216,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(196012,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(197792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(199556,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(201303,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(203033,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(204745,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(206438,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(208113,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(209769,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(211406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(213023,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(214620,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(216196,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(217751,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(219284,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(220796,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(222286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(223753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(225197,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(226619,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(228016,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(229390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(230739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(232064,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(233364,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(234638,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(235887,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(237111,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(238308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(239478,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(240622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(241739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(242828,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(243890,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(244924,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(245930,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(246908,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(247857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(248777,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(249669,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(250530,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(251363,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252166,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(253682,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(254394,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255076,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255728,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256349,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(257497,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258025,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258986,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259420,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260191,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260529,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261109,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261561,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261884,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261997,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262078,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262143,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262078,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261997,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261884,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261561,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261109,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260529,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260191,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259420,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258986,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258025,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(257497,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256349,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255728,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255076,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(254394,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(253682,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252166,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(251363,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(250530,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(249669,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(248777,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(247857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(246908,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(245930,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(244924,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(243890,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(242828,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(241739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(240622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(239478,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(238308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(237111,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(235887,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(234638,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(233364,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(232064,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(230739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(229390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(228016,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(226619,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(225197,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(223753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(222286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(220796,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(219284,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(217751,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(216196,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(214620,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(213023,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(211406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(209769,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(208113,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(206438,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(204745,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(203033,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(201303,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(199556,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(197792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(196012,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(194216,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(192404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(190577,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(188735,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(186879,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(185009,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(183126,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(181230,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(179322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(177402,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(175470,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(173528,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(171575,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(169612,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(167639,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(165658,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(163668,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(161670,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(159664,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(157651,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(155632,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(153607,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(151576,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(149540,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(147499,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(145455,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(143406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(141355,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(139302,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(137246,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(135189,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(133130,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(131072,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(129013,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(126954,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(124897,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(122841,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(120788,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(118737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(116688,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(114644,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(112603,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(110567,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(108536,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(106511,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(104492,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(102479,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(100473,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(98475,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(96485,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(94504,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(92531,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(90568,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(88615,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(86673,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(84741,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(82821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(80913,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(79017,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(77134,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(75264,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(73408,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(71566,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(69739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(67927,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(66131,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(64351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(62587,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(60840,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(59110,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(57398,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(55705,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(54030,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(52374,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(50737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(49120,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(47523,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(45947,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(44392,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(42859,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(41347,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(39857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(38390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(36946,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(35524,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(34127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(32753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(31404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(30079,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(28779,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(27505,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(26256,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(25032,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(23835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(22665,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(21521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(20404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(19315,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(18253,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(17219,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16213,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(15235,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(14286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(13366,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(12474,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(11613,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(10780,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9977,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(8461,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7749,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7067,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(6415,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5794,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4646,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4118,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3157,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2723,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1952,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1614,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1034,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(582,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(146,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(65,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(0,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(65,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(146,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(582,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1034,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1614,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1952,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2723,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3157,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4118,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4646,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5794,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(6415,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7067,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7749,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(8461,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9977,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(10780,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(11613,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(12474,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(13366,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(14286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(15235,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16213,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(17219,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(18253,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(19315,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(20404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(21521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(22665,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(23835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(25032,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(26256,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(27505,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(28779,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(30079,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(31404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(32753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(34127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(35524,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(36946,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(38390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(39857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(41347,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(42859,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(44392,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(45947,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(47523,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(49120,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(50737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(52374,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(54030,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(55705,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(57398,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(59110,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(60840,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(62587,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(64351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(66131,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(67927,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(69739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(71566,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(73408,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(75264,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(77134,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(79017,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(80913,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(82821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(84741,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(86673,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(88615,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(90568,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(92531,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(94504,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(96485,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(98475,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(100473,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(102479,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(104492,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(106511,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(108536,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(110567,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(112603,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(114644,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(116688,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(118737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(120788,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(122841,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(124897,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(126954,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(129013,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(131071,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(133130,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(135189,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(137246,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(139302,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(141355,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(143406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(145455,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(147499,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(149540,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(151576,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(153607,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(155632,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(157651,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(159664,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(161670,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(163668,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(165658,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(167639,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(169612,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(171575,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(173528,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(175470,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(177402,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(179322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(181230,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(183126,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(185009,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(186879,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(188735,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(190577,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(192404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(194216,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(196012,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(197792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(199556,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(201303,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(203033,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(204745,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(206438,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(208113,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(209769,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(211406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(213023,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(214620,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(216196,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(217751,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(219284,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(220796,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(222286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(223753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(225197,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(226619,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(228016,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(229390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(230739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(232064,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(233364,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(234638,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(235887,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(237111,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(238308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(239478,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(240622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(241739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(242828,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(243890,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(244924,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(245930,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(246908,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(247857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(248777,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(249669,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(250530,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(251363,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252166,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(253682,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(254394,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255076,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255728,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256349,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(257497,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258025,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258986,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259420,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260191,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260529,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261109,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261561,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261884,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261997,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262078,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262143,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262078,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261997,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261884,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261561,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261109,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260529,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260191,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259420,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258986,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258025,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(257497,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256349,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255728,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255076,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(254394,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(253682,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252166,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(251363,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(250530,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(249669,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(248777,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(247857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(246908,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(245930,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(244924,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(243890,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(242828,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(241739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(240622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(239478,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(238308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(237111,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(235887,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(234638,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(233364,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(232064,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(230739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(229390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(228016,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(226619,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(225197,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(223753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(222286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(220796,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(219284,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(217751,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(216196,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(214620,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(213023,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(211406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(209769,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(208113,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(206438,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(204745,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(203033,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(201303,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(199556,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(197792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(196012,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(194216,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(192404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(190577,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(188735,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(186879,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(185009,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(183126,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(181230,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(179322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(177402,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(175470,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(173528,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(171575,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(169612,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(167639,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(165658,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(163668,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(161670,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(159664,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(157651,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(155632,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(153607,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(151576,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(149540,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(147499,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(145455,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(143406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(141355,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(139302,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(137246,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(135189,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(133130,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(131072,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(129013,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(126954,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(124897,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(122841,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(120788,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(118737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(116688,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(114644,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(112603,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(110567,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(108536,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(106511,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(104492,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(102479,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(100473,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(98475,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(96485,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(94504,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(92531,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(90568,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(88615,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(86673,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(84741,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(82821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(80913,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(79017,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(77134,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(75264,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(73408,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(71566,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(69739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(67927,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(66131,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(64351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(62587,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(60840,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(59110,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(57398,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(55705,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(54030,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(52374,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(50737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(49120,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(47523,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(45947,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(44392,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(42859,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(41347,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(39857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(38390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(36946,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(35524,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(34127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(32753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(31404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(30079,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(28779,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(27505,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(26256,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(25032,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(23835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(22665,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(21521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(20404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(19315,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(18253,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(17219,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16213,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(15235,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(14286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(13366,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(12474,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(11613,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(10780,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9977,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(8461,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7749,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7067,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(6415,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5794,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4646,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4118,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3157,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2723,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1952,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1614,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1034,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(582,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(146,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(65,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(0,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(65,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(146,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(582,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1034,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1614,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1952,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2723,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3157,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4118,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4646,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5794,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(6415,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7067,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7749,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(8461,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9977,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(10780,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(11613,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(12474,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(13366,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(14286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(15235,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16213,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(17219,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(18253,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(19315,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(20404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(21521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(22665,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(23835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(25032,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(26256,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(27505,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(28779,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(30079,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(31404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(32753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(34127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(35524,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(36946,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(38390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(39857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(41347,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(42859,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(44392,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(45947,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(47523,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(49120,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(50737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(52374,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(54030,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(55705,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(57398,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(59110,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(60840,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(62587,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(64351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(66131,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(67927,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(69739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(71566,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(73408,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(75264,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(77134,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(79017,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(80913,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(82821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(84741,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(86673,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(88615,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(90568,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(92531,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(94504,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(96485,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(98475,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(100473,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(102479,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(104492,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(106511,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(108536,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(110567,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(112603,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(114644,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(116688,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(118737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(120788,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(122841,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(124897,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(126954,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(129013,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(131071,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(133130,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(135189,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(137246,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(139302,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(141355,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(143406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(145455,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(147499,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(149540,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(151576,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(153607,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(155632,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(157651,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(159664,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(161670,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(163668,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(165658,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(167639,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(169612,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(171575,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(173528,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(175470,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(177402,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(179322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(181230,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(183126,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(185009,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(186879,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(188735,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(190577,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(192404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(194216,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(196012,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(197792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(199556,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(201303,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(203033,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(204745,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(206438,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(208113,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(209769,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(211406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(213023,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(214620,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(216196,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(217751,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(219284,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(220796,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(222286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(223753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(225197,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(226619,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(228016,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(229390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(230739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(232064,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(233364,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(234638,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(235887,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(237111,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(238308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(239478,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(240622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(241739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(242828,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(243890,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(244924,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(245930,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(246908,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(247857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(248777,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(249669,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(250530,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(251363,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252166,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(253682,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(254394,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255076,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255728,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256349,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(257497,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258025,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258986,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259420,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260191,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260529,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261109,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261561,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261884,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261997,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262078,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262143,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(262078,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261997,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261884,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261561,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(261109,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260529,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(260191,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259420,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258986,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(258025,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(257497,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(256349,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255728,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(255076,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(254394,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(253682,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252939,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(252166,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(251363,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(250530,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(249669,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(248777,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(247857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(246908,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(245930,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(244924,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(243890,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(242828,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(241739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(240622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(239478,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(238308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(237111,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(235887,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(234638,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(233364,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(232064,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(230739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(229390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(228016,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(226619,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(225197,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(223753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(222286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(220796,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(219284,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(217751,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(216196,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(214620,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(213023,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(211406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(209769,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(208113,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(206438,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(204745,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(203033,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(201303,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(199556,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(197792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(196012,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(194216,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(192404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(190577,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(188735,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(186879,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(185009,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(183126,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(181230,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(179322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(177402,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(175470,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(173528,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(171575,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(169612,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(167639,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(165658,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(163668,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(161670,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(159664,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(157651,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(155632,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(153607,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(151576,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(149540,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(147499,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(145455,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(143406,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(141355,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(139302,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(137246,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(135189,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(133130,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(131071,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(129013,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(126954,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(124897,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(122841,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(120788,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(118737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(116688,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(114644,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(112603,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(110567,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(108536,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(106511,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(104492,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(102479,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(100473,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(98475,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(96485,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(94504,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(92531,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(90568,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(88615,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(86673,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(84741,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(82821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(80913,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(79017,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(77134,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(75264,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(73408,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(71566,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(69739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(67927,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(66131,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(64351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(62587,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(60840,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(59110,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(57398,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(55705,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(54030,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(52374,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(50737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(49120,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(47523,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(45947,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(44392,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(42859,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(41347,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(39857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(38390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(36946,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(35524,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(34127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(32753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(31404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(30079,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(28779,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(27505,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(26256,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(25032,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(23835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(22665,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(21521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(20404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(19315,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(18253,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(17219,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16213,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(15235,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(14286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(13366,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(12474,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(11613,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(10780,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9977,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(8461,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7749,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7067,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(6415,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5794,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4646,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4118,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3157,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2723,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1952,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1614,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1034,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(582,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(146,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(65,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(0,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(65,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(146,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(259,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(582,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(792,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1034,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1308,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1614,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(1952,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2322,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(2723,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3157,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(3622,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4118,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(4646,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(5794,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(6415,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7067,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(7749,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(8461,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9204,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(9977,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(10780,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(11613,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(12474,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(13366,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(14286,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(15235,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(16213,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(17219,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(18253,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(19315,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(20404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(21521,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(22665,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(23835,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(25032,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(26256,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(27505,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(28779,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(30079,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(31404,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(32753,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(34127,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(35524,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(36946,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(38390,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(39857,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(41347,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(42859,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(44392,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(45947,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(47523,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(49120,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(50737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(52374,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(54030,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(55705,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(57398,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(59110,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(60840,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(62587,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(64351,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(66131,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(67927,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(69739,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(71566,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(73408,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(75264,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(77134,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(79017,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(80913,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(82821,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(84741,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(86673,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(88615,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(90568,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(92531,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(94504,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(96485,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(98475,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(100473,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(102479,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(104492,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(106511,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(108536,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(110567,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(112603,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(114644,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(116688,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(118737,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(120788,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(122841,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(124897,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(126954,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);

data_i_1 <= std_logic_vector(to_unsigned(129013,18));
wait for clk_period;
write(l,to_integer(signed(data_o_4)));
writeline(f,l);


		
		
		
		
		
      -- insert stimulus here 
		file_close(f);
      wait;
   end process;

END;
